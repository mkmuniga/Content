`ifdef UVM_NO_DEPRECATED
 `define uvm_sequencer_utils(T) `uvm_component_utils(T)
`endif
